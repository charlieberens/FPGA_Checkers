module SensorManager(
    output reg [31:0] reading
)

endmodule